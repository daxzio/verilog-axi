/*

Copyright (c) 2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

//`resetall `timescale 1ns / 1ps `default_nettype none

/*
 * AXI4 config write
 */
module axi_config_wr #(
    // Width of address bus in bits
    parameter ADDR_WIDTH    = 32,
    // Width of input (slave) interface data bus in bits
    parameter DATA_WIDTH    = 32,
    // Width of input (slave) interface wstrb (width of data bus in words)
    parameter STRB_WIDTH    = (DATA_WIDTH / 8),
    // Width of ID signal
    parameter ID_WIDTH      = 8,
    // Propagate awuser signal
    parameter AWUSER_ENABLE = 0,
    // Width of awuser signal
    parameter AWUSER_WIDTH  = 1,
    // Propagate wuser signal
    parameter WUSER_ENABLE  = 0,
    // Width of wuser signal
    parameter WUSER_WIDTH   = 1,
    // Propagate buser signal
    parameter BUSER_ENABLE  = 0,
    // Width of buser signal
    parameter BUSER_WIDTH   = 1
) (
    input wire clk,
    input wire rst,

    /*
     * AXI slave interface
     */
    input  wire [    ID_WIDTH-1:0] s_axi_awid,
    input  wire [  ADDR_WIDTH-1:0] s_axi_awaddr,
    input  wire [             7:0] s_axi_awlen,
    input  wire [             2:0] s_axi_awsize,
    input  wire [             1:0] s_axi_awburst,
    input  wire                    s_axi_awlock,
    input  wire [             3:0] s_axi_awcache,
    input  wire [             2:0] s_axi_awprot,
    input  wire [             3:0] s_axi_awqos,
    input  wire [             3:0] s_axi_awregion,
    input  wire [AWUSER_WIDTH-1:0] s_axi_awuser,
    input  wire                    s_axi_awvalid,
    output wire                    s_axi_awready,
    input  wire [  DATA_WIDTH-1:0] s_axi_wdata,
    input  wire [  STRB_WIDTH-1:0] s_axi_wstrb,
    input  wire                    s_axi_wlast,
    input  wire [ WUSER_WIDTH-1:0] s_axi_wuser,
    input  wire                    s_axi_wvalid,
    output wire                    s_axi_wready,
    output wire [    ID_WIDTH-1:0] s_axi_bid,
    output wire [             1:0] s_axi_bresp,
    output wire [ BUSER_WIDTH-1:0] s_axi_buser,
    output wire                    s_axi_bvalid,
    input  wire                    s_axi_bready,

    output wire                  wr,
    output wire [ADDR_WIDTH-1:0] waddr,
    output wire [DATA_WIDTH-1:0] wdata,
    output wire [STRB_WIDTH-1:0] wstrb
);

    parameter WORD_WIDTH = STRB_WIDTH;
    parameter WORD_SIZE = DATA_WIDTH / WORD_WIDTH;

    // bus width assertions
    initial begin
        if (WORD_SIZE * STRB_WIDTH != DATA_WIDTH) begin
            $error("Error: AXI slave interface data width not evenly divisble (instance %m)");
            $finish;
        end
    end

    localparam [1:0] STATE_IDLE = 2'd0, STATE_DATA = 2'd1, STATE_DATA_2 = 2'd2, STATE_RESP = 2'd3;

    reg [1:0] state_reg = STATE_IDLE, state_next;

    reg [ID_WIDTH-1:0] id_reg = {ID_WIDTH{1'b0}}, id_next;
    reg [ADDR_WIDTH-1:0] addr_reg = {ADDR_WIDTH{1'b0}}, addr_next;
    reg [DATA_WIDTH-1:0] data_reg = {DATA_WIDTH{1'b0}}, data_next;
    reg [STRB_WIDTH-1:0] strb_reg = {STRB_WIDTH{1'b0}}, strb_next;
    reg [WUSER_WIDTH-1:0] wuser_reg = {WUSER_WIDTH{1'b0}}, wuser_next;
    reg [ADDR_WIDTH-1:0] waddr_reg = {ADDR_WIDTH{1'b0}}, waddr_next;
    reg wr_reg = 1'b0, wr_next;

    reg s_axi_awready_reg = 1'b0, s_axi_awready_next;
    reg s_axi_wready_reg = 1'b0, s_axi_wready_next;
    reg [ID_WIDTH-1:0] s_axi_bid_reg = {ID_WIDTH{1'b0}}, s_axi_bid_next;
    reg [1:0] s_axi_bresp_reg = 2'd0, s_axi_bresp_next;
    reg [BUSER_WIDTH-1:0] s_axi_buser_reg = {BUSER_WIDTH{1'b0}}, s_axi_buser_next;
    reg s_axi_bvalid_reg = 1'b0, s_axi_bvalid_next;

    assign s_axi_awready = s_axi_awready_reg;
    assign s_axi_wready  = s_axi_wready_reg;
    assign s_axi_bid     = s_axi_bid_reg;
    assign s_axi_bresp   = s_axi_bresp_reg;
    assign s_axi_buser   = BUSER_ENABLE ? s_axi_buser_reg : {BUSER_WIDTH{1'b0}};
    assign s_axi_bvalid  = s_axi_bvalid_reg;

    assign waddr         = waddr_reg;
    assign wdata         = data_reg;
    assign wstrb         = strb_reg;
    assign wr            = wr_reg;

    always @(*) begin
        state_next         = STATE_IDLE;

        id_next            = id_reg;
        addr_next          = addr_reg;
        data_next          = data_reg;
        strb_next          = strb_reg;
        wuser_next         = wuser_reg;

        s_axi_awready_next = 1'b0;
        s_axi_wready_next  = 1'b0;
        s_axi_bid_next     = s_axi_bid_reg;
        s_axi_bresp_next   = s_axi_bresp_reg;
        s_axi_buser_next   = s_axi_buser_reg;
        s_axi_bvalid_next  = s_axi_bvalid_reg && !s_axi_bready;

        waddr_next = waddr_reg;
        wr_next    = 0;


        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                //s_axi_awready_next = !m_axi_awvalid;
                s_axi_awready_next = 1;

                addr_next = s_axi_awaddr;
                if (s_axi_awready && s_axi_awvalid) begin
                    s_axi_awready_next = 1'b0;
                    id_next            = s_axi_awid;
                    strb_next          = s_axi_wstrb;
                    state_next         = STATE_DATA;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                // data state; transfer write data
                s_axi_wready_next = 1;

//                 if (s_axi_wready && s_axi_wvalid) begin
//                 end
                if (s_axi_wready && s_axi_wvalid) begin
                    addr_next  = addr_reg + 4;
                    waddr_next = addr_reg;
                    wr_next    = 1;
                    data_next  = s_axi_wdata;
                    if (s_axi_wlast) begin
                        // last data word, wait for response
                        s_axi_wready_next = 1'b0;
                        state_next        = STATE_RESP;
                    end else begin
                        state_next = STATE_DATA;
                    end
                end else begin
                    state_next = STATE_DATA;
                end
            end
            STATE_RESP: begin
                // resp state; transfer write response
                s_axi_bid_next     = id_reg;
                s_axi_bresp_next   = 0;
                s_axi_buser_next   = 0;
                s_axi_bvalid_next  = 1'b1;
                s_axi_awready_next = 1;
                state_next         = STATE_IDLE;
            end
            default: state_next    = STATE_IDLE;
        endcase
    end

    always @(posedge clk) begin
        state_reg         <= state_next;

        id_reg            <= id_next;
        addr_reg          <= addr_next;
        data_reg          <= data_next;
        strb_reg          <= strb_next;
        wuser_reg         <= wuser_next;
        waddr_reg         <= waddr_next;
        wr_reg            <= wr_next;

        s_axi_awready_reg <= s_axi_awready_next;
        s_axi_wready_reg  <= s_axi_wready_next;
        s_axi_bid_reg     <= s_axi_bid_next;
        s_axi_bresp_reg   <= s_axi_bresp_next;
        s_axi_buser_reg   <= s_axi_buser_next;
        s_axi_bvalid_reg  <= s_axi_bvalid_next;

        if (rst) begin
            state_reg         <= STATE_IDLE;

            s_axi_awready_reg <= 1'b0;
            s_axi_wready_reg  <= 1'b0;
            s_axi_bvalid_reg  <= 1'b0;

        end
    end

endmodule

`resetall
